module debounce_count(input button, input reset, clk, outleds);
	output [7:0] outleds;
	reg [7:0] answer;
	reg  button_reg;
	reg  button_sync;
	wire button_done;
	wire button_click;
	reg [7:0] button_count;
	reg [7:0] outleds;

	parameter DEBOUNCE_DELAY = 32'd0_500_000;   /// 10nS * 1M = 10mS

	always @(posedge clk)   button_reg   <= button;
	always @(posedge clk)   button_sync  <= !button_reg;

	assign	button_done  = (button_count == DEBOUNCE_DELAY); 
	assign	button_click = (button_count == DEBOUNCE_DELAY - 1); 

	always @(posedge clk) 
        	  if (!button_sync)      button_count <= 0;
          	else if (button_done)  button_count <= button_count;
          	else                   button_count <= button_count + 1;

	always @(posedge clk)
		if (button_click)	answer <= answer + 1;
		else if (!reset)	answer <= 0;
		else			answer <= answer;
		
	always @(answer)
		case(cathode_select)
			0: outleds <= 8'b0000_0000;
			1: outleds <= 8'b0000_0000;
			2: outleds <= 8'b0000_0000;
			3: outleds <= 8'b0000_0000;
			4: outleds <= 8'b0000_0000;
			5: outleds <= 8'b0000_0000;
endmodule
