`timescale 1ns / 1ps

module State(sw1, sw2, button, detected_signal);
input sw1;
input sw2;
input button;
output detected signal;


endmodule
